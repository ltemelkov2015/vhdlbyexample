-- This is the whole module that talk to USB MCU